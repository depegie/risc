`ifndef DEFINES_VH
`define DEFINES_VH

`define RAM_CAPACITY 'd16
`define WORD_SIZE 'd4

`endif