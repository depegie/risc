module uart_tx (
    input         Clk,
    input         Rst,
    output        Tx,
    input [7 : 0] S_axis_tdata,
    input         S_axis_tvalid,
    output        S_axis_tready
);


endmodule