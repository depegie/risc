interface monitor_if;
    logic rx;
endinterface