interface driver_if;
    logic tx;
endinterface