`ifndef DEFINES_VH
`define DEFINES_VH

`define RAM_CAPACITY  'd128
`define ADDR_SIZE     $clog2(`RAM_CAPACITY)
`define WORD_SIZE_B   'd4

`endif