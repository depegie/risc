`ifndef DEFINES_SVH
`define DEFINES_SVH

`define RAM_CAPACITY_B 128
`define ADDR_SIZE      $clog2(`RAM_CAPACITY_B)
`define WORD_SIZE_B    4
`define WORD_SIZE      8*`WORD_SIZE_B

`endif